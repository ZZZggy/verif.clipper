//------------------------------------------------------------------------------
// ACCEDIAN NETWORKS
// High Performance Service Assurance (TM)
//
// Accedian Networks, Inc.
// 4878 Levy, suite 202
// Saint-Laurent, Quebec Canada H4R 2P1
// E-mail: support@accedian.com
// Website: www.accedian.com
//
// ACCEDIAN PROPRIETARY
//
// COPYRIGHT (c) BY ACCEDIAN CORPORATION. ALL RIGHTS RESERVED. NO
// PART OF THIS PROGRAM OR PUBLICATION MAY BE REPRODUCED, TRANSMITTED,
// TRANSCRIBED, STORED IN A RETRIEVAL SYSTEM, OR TRANSLATED INTO ANY LANGUAGE
// OR COMPUTER LANGUAGE IN ANY FORM OR BY ANY MEANS, ELECTRONIC, MECHANICAL,
// MAGNETIC, OPTICAL, CHEMICAL, MANUAL, OR OTHERWISE, WITHOUT THE PRIOR
// WRITTEN PERMISSION OF ACCEDIAN INC.
//
//------------------------------------------------------------------------------
// !!! AUTO-GENERATED FILE !!!
// Register definitions for altera_xcvr_reconfig register block.
//
// To enable per-instance coverage: regmodel...set_per_instance_coverage(1, UVM_(NO_)HIER);
// To enable singleton coverage:    regmodel...set_per_instance_coverage(0, UVM_(NO_)HIER);
// To enable coverage:              void'(regmodel...set_coverage(1));
// To enable hierarchical coverage: void'(regmodel...set_coverage(UVM_CVR_ALL));
//
// TODO: <field>.configure: need to replace:has_reset => actual, individually_accessible => byte lane accessible
// TODO: add address coverage to register blocks
// TODO: for memories in blocks, n_bits and access should be configured somehow
//       mem = new("mem", addressRange, `UVM_REG_DATA_WIDTH, "RW", UVM_NO_COVERAGE); // mem_type::type_id::create("mem", , get_full_name());
// TODO: for block default_map, specify actual n_bytes, endian-ness, byte_addressing
//------------------------------------------------------------------------------

`include "uvm_macros.svh"

//---------------------------------------------------------
// Group: altera_xcvr_reconfig
//---------------------------------------------------------

package altera_xcvr_reconfig_reg_pkg;
    import uvm_pkg::*;
    import acd_uvm_pkg::*;
    import pma_analog_control_regiters_reg_pkg::*;
    import atx_pll_cal_registers_reg_pkg::*;
    import streamer_module_registers_reg_pkg::*;
    import pll_reconfiguration_registers_reg_pkg::*;
    import dcd_calibration_registers_reg_pkg::*;






// Class: altera_xcvr_reconfig_reg_block
// Register Block .altera_xcvr_reconfig: 
class altera_xcvr_reconfig_reg_block extends uvm_reg_block;

    // Validate register width
    local static bit valid_reg_data_width = check_data_width(`UVM_REG_DATA_WIDTH);

    rand pma_analog_control_regiters_reg_block pma_analog_control_regiters;
    rand atx_pll_cal_registers_reg_block atx_pll_cal_registers;
    rand streamer_module_registers_reg_block streamer_module_registers;
    rand pll_reconfiguration_registers_reg_block pll_reconfiguration_registers;
    rand dcd_calibration_registers_reg_block dcd_calibration_registers;

    // Variable: params
    // Parameter key/value lookup.
    static protected acd_reg_param_cfg m_params;

    // Variable: cg_per_instance
    // Assert to construct all sub-block and register covergroups per instance rather than singleton
    protected bit cg_per_instance;

    `uvm_object_utils(altera_xcvr_reconfig_reg_pkg::altera_xcvr_reconfig_reg_block)

    // Constructor: new
    function new(string name = "altera_xcvr_reconfig_reg_block");
        super.new(name, UVM_NO_COVERAGE);
    endfunction


    // Function: build
    virtual function void build();
        if ((m_params == null) && (0 > 0))
            if (!uvm_config_db#(acd_reg_param_cfg)::get(null, get_full_name(), "cfg", m_params))
                `uvm_fatal("CFGERR", {get_full_name(), " failed to get configuration for parameters."})


        pma_analog_control_regiters = pma_analog_control_regiters_reg_block::type_id::create("pma_analog_control_regiters", , get_full_name());
        atx_pll_cal_registers = atx_pll_cal_registers_reg_block::type_id::create("atx_pll_cal_registers", , get_full_name());
        streamer_module_registers = streamer_module_registers_reg_block::type_id::create("streamer_module_registers", , get_full_name());
        pll_reconfiguration_registers = pll_reconfiguration_registers_reg_block::type_id::create("pll_reconfiguration_registers", , get_full_name());
        dcd_calibration_registers = dcd_calibration_registers_reg_block::type_id::create("dcd_calibration_registers", , get_full_name());

        pma_analog_control_regiters.configure(this);
        atx_pll_cal_registers.configure(this);
        streamer_module_registers.configure(this);
        pll_reconfiguration_registers.configure(this);
        dcd_calibration_registers.configure(this);

        pma_analog_control_regiters.build();
        atx_pll_cal_registers.build();
        streamer_module_registers.build();
        pll_reconfiguration_registers.build();
        dcd_calibration_registers.build();

        // define default map
        default_map = create_map("altera_xcvr_reconfig_default_map", 'h0, `UVM_REG_DATA_WIDTH/8, UVM_NO_ENDIAN, 0);
        this.default_map.add_submap(this.pma_analog_control_regiters.default_map, 'h0);
        this.default_map.add_submap(this.atx_pll_cal_registers.default_map, 'h0);
        this.default_map.add_submap(this.streamer_module_registers.default_map, 'h0);
        this.default_map.add_submap(this.pll_reconfiguration_registers.default_map, 'h0);
        this.default_map.add_submap(this.dcd_calibration_registers.default_map, 'h0);

        // Recursively lock register model and build the address map to enable
        // uvm_reg_map::get_reg_by_offset() and uvm_reg_map::get_mem_by_offset() methods.
        // It is impossible to unlock a model.
        lock_model();
    endfunction


     // Function: set_per_instance_coverage
     // Enable or disable instance coverage, otherwise singleton coverage.
     virtual function void set_per_instance_coverage(bit per_inst, uvm_hier_e hier=UVM_HIER);
         this.cg_per_instance = per_inst;

        // Use UVM_CVR_ALL for hierarchical enabling.
        if(hier == UVM_HIER) begin
            pma_analog_control_regiters.set_per_instance_coverage(per_inst, hier);
            atx_pll_cal_registers.set_per_instance_coverage(per_inst, hier);
            streamer_module_registers.set_per_instance_coverage(per_inst, hier);
            pll_reconfiguration_registers.set_per_instance_coverage(per_inst, hier);
            dcd_calibration_registers.set_per_instance_coverage(per_inst, hier);
        end
     endfunction


    // Function: set_coverage
    // Override base function to create covergroups for all registers in this block.
    //
    // In order to enable hierarchical creation, use UVM_CVR_ALL.
    virtual function uvm_reg_cvr_t set_coverage(uvm_reg_cvr_t is_on);
        //void'(uvm_config_db#(bit)::get(null, get_full_name(), "cg_per_instance", cg_per_instance));
        set_coverage = super.set_coverage(is_on);
        // Use UVM_CVR_ALL for hierarchical enabling.
        if(is_on == UVM_CVR_ALL) begin
            //void'(uvm_config_db#(bit)::set(null, pma_analog_control_regiters.get_full_name(), "cg_per_instance", cg_per_instance));
            void'(pma_analog_control_regiters.set_coverage(is_on));
            //void'(uvm_config_db#(bit)::set(null, atx_pll_cal_registers.get_full_name(), "cg_per_instance", cg_per_instance));
            void'(atx_pll_cal_registers.set_coverage(is_on));
            //void'(uvm_config_db#(bit)::set(null, streamer_module_registers.get_full_name(), "cg_per_instance", cg_per_instance));
            void'(streamer_module_registers.set_coverage(is_on));
            //void'(uvm_config_db#(bit)::set(null, pll_reconfiguration_registers.get_full_name(), "cg_per_instance", cg_per_instance));
            void'(pll_reconfiguration_registers.set_coverage(is_on));
            //void'(uvm_config_db#(bit)::set(null, dcd_calibration_registers.get_full_name(), "cg_per_instance", cg_per_instance));
            void'(dcd_calibration_registers.set_coverage(is_on));
        end
        return set_coverage;
    endfunction


    // Function: fields2string
    // Stringify.
    virtual function string convert2string();
        string s = "";
        uvm_reg regs[$];
        uvm_reg_field fields[$];

        get_registers(regs, UVM_HIER);
        $swrite(s, "\nUVM_REG_BLOCK::%0s (%0d registers)\n", get_name, regs.size());
        foreach (regs[m]) begin
            $swrite(s, "%0s    %0s=0x%16h\n", s, regs[m].get_full_name, regs[m].get());
            // Getting the fields is optional might be too verbose
            //fields.delete();
            //regs[m].get_fields(fields);
            //foreach (fields[n]) begin
                //$swrite(s, "%0s        %0s=0x%0h\n", s, fields[n].get_full_name, fields[n].value);
            //end
        end
        return s;
    endfunction


    // Function: regs2update
    // Stringifying only regmodel registers that need updating. Useful after randomization.
    virtual function string regs2update();
        string s = "";
        uvm_reg regs[$];
        uvm_reg_field fields[$];

        get_registers(regs, UVM_HIER);
        $swrite(s, "\nRegisters requiring update in UVM_REG_BLOCK::%0s\n", get_name);
        foreach (regs[m]) begin
            if (regs[m].needs_update()) begin
                $swrite(s, "%0s    %0s=0x%16h\n", s, regs[m].get_full_name, regs[m].get());
                // Getting the fields is optional might be too verbose
                fields.delete();
                regs[m].get_fields(fields);
                foreach (fields[n]) begin
                    $swrite(s, "%0s        %0s=0x%0h\n", s, fields[n].get_full_name, fields[n].value);
                end
            end
        end
        return s;
    endfunction

endclass

endpackage