//------------------------------------------------------------------------------
// ACCEDIAN NETWORKS
// High Performance Service Assurance (TM)
//
// Accedian Networks, Inc.
// 4878 Levy, suite 202
// Saint-Laurent, Quebec Canada H4R 2P1
// E-mail: support@accedian.com
// Website: www.accedian.com
//
// ACCEDIAN PROPRIETARY
//
// COPYRIGHT (c) BY ACCEDIAN CORPORATION. ALL RIGHTS RESERVED. NO
// PART OF THIS PROGRAM OR PUBLICATION MAY BE REPRODUCED, TRANSMITTED,
// TRANSCRIBED, STORED IN A RETRIEVAL SYSTEM, OR TRANSLATED INTO ANY LANGUAGE
// OR COMPUTER LANGUAGE IN ANY FORM OR BY ANY MEANS, ELECTRONIC, MECHANICAL,
// MAGNETIC, OPTICAL, CHEMICAL, MANUAL, OR OTHERWISE, WITHOUT THE PRIOR
// WRITTEN PERMISSION OF ACCEDIAN INC.
//
//------------------------------------------------------------------------------
// !!! AUTO-GENERATED FILE !!!
// Register definitions for mac10g_if register block.
//
// To enable per-instance coverage: regmodel...set_per_instance_coverage(1, UVM_(NO_)HIER);
// To enable singleton coverage:    regmodel...set_per_instance_coverage(0, UVM_(NO_)HIER);
// To enable coverage:              void'(regmodel...set_coverage(1));
// To enable hierarchical coverage: void'(regmodel...set_coverage(UVM_CVR_ALL));
//
// TODO: <field>.configure: need to replace:has_reset => actual, individually_accessible => byte lane accessible
// TODO: add address coverage to register blocks
// TODO: for memories in blocks, n_bits and access should be configured somehow
//       mem = new("mem", addressRange, `UVM_REG_DATA_WIDTH, "RW", UVM_NO_COVERAGE); // mem_type::type_id::create("mem", , get_full_name());
// TODO: for block default_map, specify actual n_bytes, endian-ness, byte_addressing
//------------------------------------------------------------------------------

`include "uvm_macros.svh"

//---------------------------------------------------------
// Group: mac10g_if
//---------------------------------------------------------

package mac10g_if_reg_pkg;
    import uvm_pkg::*;
    import acd_uvm_pkg::*;
    import xgmac_rx_cfg_reg_pkg::*;
    import xgmac_rx_stats_reg_pkg::*;
    import xgmac_tx_cfg_reg_pkg::*;
    import xgmac_tx_stats_reg_pkg::*;






// Class: mac10g_if_reg_block
// Register Block .mac10g_if: 
class mac10g_if_reg_block extends uvm_reg_block;

    // Validate register width
    local static bit valid_reg_data_width = check_data_width(`UVM_REG_DATA_WIDTH);

    rand xgmac_rx_cfg_reg_block xgmac_rx_cfg;
    rand xgmac_rx_stats_reg_block xgmac_rx_stats;
    rand xgmac_tx_cfg_reg_block xgmac_tx_cfg;
    rand xgmac_tx_stats_reg_block xgmac_tx_stats;

    // Variable: params
    // Parameter key/value lookup.
    static protected acd_reg_param_cfg m_params;

    // Variable: cg_per_instance
    // Assert to construct all sub-block and register covergroups per instance rather than singleton
    protected bit cg_per_instance;

    `uvm_object_utils(mac10g_if_reg_pkg::mac10g_if_reg_block)

    // Constructor: new
    function new(string name = "mac10g_if_reg_block");
        super.new(name, UVM_NO_COVERAGE);
    endfunction


    // Function: build
    virtual function void build();
        if ((m_params == null) && (0 > 0))
            if (!uvm_config_db#(acd_reg_param_cfg)::get(null, get_full_name(), "cfg", m_params))
                `uvm_fatal("CFGERR", {get_full_name(), " failed to get configuration for parameters."})


        xgmac_rx_cfg = xgmac_rx_cfg_reg_block::type_id::create("xgmac_rx_cfg", , get_full_name());
        xgmac_rx_stats = xgmac_rx_stats_reg_block::type_id::create("xgmac_rx_stats", , get_full_name());
        xgmac_tx_cfg = xgmac_tx_cfg_reg_block::type_id::create("xgmac_tx_cfg", , get_full_name());
        xgmac_tx_stats = xgmac_tx_stats_reg_block::type_id::create("xgmac_tx_stats", , get_full_name());

        xgmac_rx_cfg.configure(this);
        xgmac_rx_stats.configure(this);
        xgmac_tx_cfg.configure(this);
        xgmac_tx_stats.configure(this);

        xgmac_rx_cfg.build();
        xgmac_rx_stats.build();
        xgmac_tx_cfg.build();
        xgmac_tx_stats.build();

        // define default map
        default_map = create_map("mac10g_if_default_map", 'h0, `UVM_REG_DATA_WIDTH/8, UVM_NO_ENDIAN, 0);
        this.default_map.add_submap(this.xgmac_rx_cfg.default_map, 'h0);
        this.default_map.add_submap(this.xgmac_rx_stats.default_map, 'h80);
        this.default_map.add_submap(this.xgmac_tx_cfg.default_map, 'h100);
        this.default_map.add_submap(this.xgmac_tx_stats.default_map, 'h180);

        // Recursively lock register model and build the address map to enable
        // uvm_reg_map::get_reg_by_offset() and uvm_reg_map::get_mem_by_offset() methods.
        // It is impossible to unlock a model.
        lock_model();
    endfunction


     // Function: set_per_instance_coverage
     // Enable or disable instance coverage, otherwise singleton coverage.
     virtual function void set_per_instance_coverage(bit per_inst, uvm_hier_e hier=UVM_HIER);
         this.cg_per_instance = per_inst;

        // Use UVM_CVR_ALL for hierarchical enabling.
        if(hier == UVM_HIER) begin
            xgmac_rx_cfg.set_per_instance_coverage(per_inst, hier);
            xgmac_rx_stats.set_per_instance_coverage(per_inst, hier);
            xgmac_tx_cfg.set_per_instance_coverage(per_inst, hier);
            xgmac_tx_stats.set_per_instance_coverage(per_inst, hier);
        end
     endfunction


    // Function: set_coverage
    // Override base function to create covergroups for all registers in this block.
    //
    // In order to enable hierarchical creation, use UVM_CVR_ALL.
    virtual function uvm_reg_cvr_t set_coverage(uvm_reg_cvr_t is_on);
        //void'(uvm_config_db#(bit)::get(null, get_full_name(), "cg_per_instance", cg_per_instance));
        set_coverage = super.set_coverage(is_on);
        // Use UVM_CVR_ALL for hierarchical enabling.
        if(is_on == UVM_CVR_ALL) begin
            //void'(uvm_config_db#(bit)::set(null, xgmac_rx_cfg.get_full_name(), "cg_per_instance", cg_per_instance));
            void'(xgmac_rx_cfg.set_coverage(is_on));
            //void'(uvm_config_db#(bit)::set(null, xgmac_rx_stats.get_full_name(), "cg_per_instance", cg_per_instance));
            void'(xgmac_rx_stats.set_coverage(is_on));
            //void'(uvm_config_db#(bit)::set(null, xgmac_tx_cfg.get_full_name(), "cg_per_instance", cg_per_instance));
            void'(xgmac_tx_cfg.set_coverage(is_on));
            //void'(uvm_config_db#(bit)::set(null, xgmac_tx_stats.get_full_name(), "cg_per_instance", cg_per_instance));
            void'(xgmac_tx_stats.set_coverage(is_on));
        end
        return set_coverage;
    endfunction


    // Function: fields2string
    // Stringify.
    virtual function string convert2string();
        string s = "";
        uvm_reg regs[$];
        uvm_reg_field fields[$];

        get_registers(regs, UVM_HIER);
        $swrite(s, "\nUVM_REG_BLOCK::%0s (%0d registers)\n", get_name, regs.size());
        foreach (regs[m]) begin
            $swrite(s, "%0s    %0s=0x%16h\n", s, regs[m].get_full_name, regs[m].get());
            // Getting the fields is optional might be too verbose
            //fields.delete();
            //regs[m].get_fields(fields);
            //foreach (fields[n]) begin
                //$swrite(s, "%0s        %0s=0x%0h\n", s, fields[n].get_full_name, fields[n].value);
            //end
        end
        return s;
    endfunction


    // Function: regs2update
    // Stringifying only regmodel registers that need updating. Useful after randomization.
    virtual function string regs2update();
        string s = "";
        uvm_reg regs[$];
        uvm_reg_field fields[$];

        get_registers(regs, UVM_HIER);
        $swrite(s, "\nRegisters requiring update in UVM_REG_BLOCK::%0s\n", get_name);
        foreach (regs[m]) begin
            if (regs[m].needs_update()) begin
                $swrite(s, "%0s    %0s=0x%16h\n", s, regs[m].get_full_name, regs[m].get());
                // Getting the fields is optional might be too verbose
                fields.delete();
                regs[m].get_fields(fields);
                foreach (fields[n]) begin
                    $swrite(s, "%0s        %0s=0x%0h\n", s, fields[n].get_full_name, fields[n].value);
                end
            end
        end
        return s;
    endfunction

endclass

endpackage