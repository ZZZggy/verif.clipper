`include "shaper_group_1_regs.svh"
`include "shaper_group_0_regs.svh"
`include "uni_q_stats_regs.svh"
`include "nni1_q_stats_regs.svh"
`include "nni0_q_stats_regs.svh"
`include "uni_q_system_regs.svh"
`include "nni1_q_system_regs.svh"
`include "nni0_q_system_regs.svh"
`include "tm_globals_regs.svh"
`include "scheduler_regs.svh"
`include "shaper_regs.svh"
`include "q_stats_regs.svh"
`include "q_system_regs.svh"
`include "cos_actions_regs.svh"
`include "cos_actions_uni1g_regs.svh"
`include "cos_actions_uni10g_regs.svh"
`include "cos_actions_nni10g_regs.svh"
`include "rule_action_mapping_uni1g_regs.svh"
`include "rule_action_mapping_uni10g_regs.svh"
`include "rule_action_mapping_nni10g_regs.svh"
`include "cos_pattern_uni1g_regs.svh"
`include "cos_pattern_uni10g_regs.svh"
`include "cos_pattern_nni10g_regs.svh"
`include "vid_table_uni1g_regs.svh"
`include "vid_table_uni10g_regs.svh"
`include "vid_table_nni10g_regs.svh"
`include "class_stats_1g_regs.svh"
`include "class_stats_10g1g_regs.svh"
`include "class_stats_10g_regs.svh"
`include "class_stats_cpu_regs.svh"
`include "class_stats_if_regs.svh"
`include "vid_pairing_table_uni1g_regs.svh"
`include "vid_pairing_table_uni10g_regs.svh"
`include "vid_pairing_table_nni10g_regs.svh"
`include "fwd_instance_memory_regs.svh"
`include "fwd_domain_memory_regs.svh"
`include "fwd_vid_memory_regs.svh"
`include "class2bwp_profile_ndx_regs.svh"
`include "profile_ndx_regs.svh"
`include "profile_cfg_ndx_regs.svh"
`include "bwp_shaper_regs.svh"
`include "bwp_profile_remap_regs.svh"
`include "bwp_profile_stats_regs.svh"
`include "bwp_profile_cfgs_regs.svh"
`include "pktgen_shapping_regs.svh"
`include "pktgen_padding_regs.svh"
`include "pktgen_flowheader_regs.svh"
`include "q_map_tbl_cos_internal_regs.svh"
`include "q_map_tbl_outgoing_qset_regs.svh"
`include "q_map_tbl_outgoing_port_regs.svh"
`include "dcd_calibration_registers_regs.svh"
`include "pll_reconfiguration_registers_regs.svh"
`include "streamer_module_registers_regs.svh"
`include "atx_pll_cal_registers_regs.svh"
`include "pma_analog_control_regiters_regs.svh"
`include "gmii_pcs_registers_regs.svh"
`include "pcs_registers_regs.svh"
`include "pma_registers_regs.svh"
`include "pcs_registers_1g_regs.svh"
`include "phy_if_globals_regs.svh"
`include "altera_xcvr_reconfig_regs.svh"
`include "altera_phy_1g10g_regs.svh"
`include "altera_phy_1g_regs.svh"
`include "xgmac_tx_stats_regs.svh"
`include "xgmac_tx_cfg_regs.svh"
`include "xgmac_rx_stats_regs.svh"
`include "xgmac_rx_cfg_regs.svh"
`include "tse_mac_stats_tx_regs.svh"
`include "tse_mac_stats_rx_regs.svh"
`include "tse_mac_tx_regs.svh"
`include "tse_mac_rx_regs.svh"
`include "tse_mac_stats_regs.svh"
`include "tse_mac_regs.svh"
`include "cos_mark_tbl_cfi_pcp_regs.svh"
`include "cos_mark_tbl_port_regs.svh"
`include "timebase2_core_compensations_regs.svh"
`include "timebase2_core_globals_regs.svh"
`include "protection_tbl_physical_port_regs.svh"
`include "protection_tbl_logical_port_regs.svh"
`include "port_input_cfg_regs.svh"
`include "access_logger_regs.svh"
`include "classifiers_regs.svh"
`include "traffic_manager_regs.svh"
`include "cpu_monitor_domain_action_regs.svh"
`include "cos_action_top_regs.svh"
`include "rule_action_mapping_top_regs.svh"
`include "cos_pattern_tables_top_regs.svh"
`include "vid_table_regs.svh"
`include "class_stats_top_regs.svh"
`include "vid_pairing_table_regs.svh"
`include "fwd_db_regs.svh"
`include "bwp_regs.svh"
`include "pktgen_regs.svh"
`include "q_map_tbl_regs.svh"
`include "phy_if_regs.svh"
`include "inspector_regs.svh"
`include "mac10g_if_regs.svh"
`include "mac_if_regs.svh"
`include "acd_seq_checker_reg_regs.svh"
`include "cos_mark_tbl_regs.svh"
`include "mem_ctrl_regs.svh"
`include "clock_ctrl_regs.svh"
`include "platform_ctrl_regs.svh"
`include "i2c_regs.svh"
`include "flush_stat_regs.svh"
`include "cpu_bucket_regs.svh"
`include "timebase2_regs.svh"
`include "protection_tbl_regs.svh"
`include "chip_global_regs.svh"
`include "c1lt_regs.svh"
