//------------------------------------------------------------------------------
// ACCEDIAN NETWORKS
// High Performance Service Assurance (TM)
//
// Accedian Networks, Inc.
// 4878 Levy, suite 202
// Saint-Laurent, Quebec Canada H4R 2P1
// E-mail: support@accedian.com
// Website: www.accedian.com
//
// ACCEDIAN PROPRIETARY
//
// COPYRIGHT (c) BY ACCEDIAN CORPORATION. ALL RIGHTS RESERVED. NO
// PART OF THIS PROGRAM OR PUBLICATION MAY BE REPRODUCED, TRANSMITTED,
// TRANSCRIBED, STORED IN A RETRIEVAL SYSTEM, OR TRANSLATED INTO ANY LANGUAGE
// OR COMPUTER LANGUAGE IN ANY FORM OR BY ANY MEANS, ELECTRONIC, MECHANICAL,
// MAGNETIC, OPTICAL, CHEMICAL, MANUAL, OR OTHERWISE, WITHOUT THE PRIOR
// WRITTEN PERMISSION OF ACCEDIAN INC.
//
//------------------------------------------------------------------------------
// !!! AUTO-GENERATED FILE !!!
// Register definitions for rule_action_mapping_nni10g register block.
//
// To enable per-instance coverage: regmodel...set_per_instance_coverage(1, UVM_(NO_)HIER);
// To enable singleton coverage:    regmodel...set_per_instance_coverage(0, UVM_(NO_)HIER);
// To enable coverage:              void'(regmodel...set_coverage(1));
// To enable hierarchical coverage: void'(regmodel...set_coverage(UVM_CVR_ALL));
//
// TODO: <field>.configure: need to replace:has_reset => actual, individually_accessible => byte lane accessible
// TODO: add address coverage to register blocks
// TODO: for memories in blocks, n_bits and access should be configured somehow
//       mem = new("mem", addressRange, `UVM_REG_DATA_WIDTH, "RW", UVM_NO_COVERAGE); // mem_type::type_id::create("mem", , get_full_name());
// TODO: for block default_map, specify actual n_bytes, endian-ness, byte_addressing
//------------------------------------------------------------------------------

`include "uvm_macros.svh"

//---------------------------------------------------------
// Group: rule_action_mapping_nni10g
//---------------------------------------------------------

package rule_action_mapping_nni10g_reg_pkg;
    import uvm_pkg::*;
    import acd_uvm_pkg::*;

typedef class p5_priority_index_reg_cover;

// Class: p5_priority_index_reg
// Register p5.priority_index: Maps the rule priority indexes from vid_table and classifiers to rule action indexes toward cos_action.
class p5_priority_index_reg extends uvm_reg;

    // Variable: if_action_index
    // remapping of if rule priority index to if_rule_action_index
    rand uvm_reg_field if_action_index;
    // Variable: cpu_action_index
    // remapping of cpu rule priority index to cpu_rule_action_index
    rand uvm_reg_field cpu_action_index;
    // Variable: mon1_action_index
    // remapping of mon1 rule priority index to mon1_rule_action_index
    rand uvm_reg_field mon1_action_index;
    // Variable: mon2_action_index
    // remapping of mon2 rule priority index to mon2_rule_action_index
    rand uvm_reg_field mon2_action_index;

    // Variable: m_params
    // Parameter key/value lookup.
    static protected acd_reg_param_cfg m_params;

    // Variable: cg
    // Coverage object. Static to reduce memory usage.
    static p5_priority_index_reg_cover cg_all;

    // Variable: cg
    // Coverage object.
    p5_priority_index_reg_cover cg;

    // Variable: is_read
    // Last access type.
    protected bit is_read;

    `uvm_object_utils(rule_action_mapping_nni10g_reg_pkg::p5_priority_index_reg)

    // Constructor: new
    function new(string name = "p5_priority_index");
        super.new(name, `UVM_REG_DATA_WIDTH, UVM_NO_COVERAGE);
    endfunction


    // Function: build
    virtual function void build();
        if ((m_params == null) && has_params())
            if (!uvm_config_db#(acd_reg_param_cfg)::get(null, get_full_name(), "cfg", m_params))
                `uvm_fatal("CFGERR", {get_full_name(), " failed to get configuration for parameters."})

        if_action_index = uvm_reg_field::type_id::create("if_action_index", , get_full_name());
        cpu_action_index = uvm_reg_field::type_id::create("cpu_action_index", , get_full_name());
        mon1_action_index = uvm_reg_field::type_id::create("mon1_action_index", , get_full_name());
        mon2_action_index = uvm_reg_field::type_id::create("mon2_action_index", , get_full_name());

        // uvm_reg_field::configure(uvm_reg parent, int unsigned size, int unsigned lsb_pos, string access, bit volatile, uvm_reg_data_t reset, bit has_reset, bit is_rand, bit individually_accessible)
        if_action_index.configure(this, 11, 0, "RW", 0, 'h0, 1, 1, 0);
        cpu_action_index.configure(this, 6, 14, "RW", 0, 'h0, 1, 1, 0);
        mon1_action_index.configure(this, 1, 24, "RW", 0, 'h0, 1, 1, 0);
        mon2_action_index.configure(this, 1, 28, "RW", 0, 'h0, 1, 1, 0);
    endfunction


    // Function: RMW
    // Helper task for read-modify-write based on mask.
    // Ones in the mask position indicate bits to modify.
    task RMW(output uvm_status_e status, input uvm_reg_data_t data, input uvm_reg_data_t mask);
        uvm_reg_data_t tmp;

        // read
        read(status, tmp);
        // modify
        tmp &= ~mask;
        tmp |= data & mask;
        //write
        write(status, tmp);
    endtask


    // Function: post_write
    // Add message after access.
    virtual task post_write(uvm_reg_item rw);
        super.post_write(rw);
        is_read = 0;
        `uvm_info("REG", $sformatf("%0s WRITE=0x%0h ADDR=0x%0h%0s", this.get_full_name(), this.get(), this.get_address(), this.fields2string()), UVM_MEDIUM)
        sample_values();
    endtask


    // Function: post_read
    // Add message after access.
    virtual task post_read(uvm_reg_item rw);
        super.post_read(rw);
        is_read = 1;
        `uvm_info("REG", $sformatf("%0s READ=0x%0h ADDR=0x%0h%0s", this.get_full_name(), this.get(), this.get_address(), this.fields2string()), UVM_MEDIUM)
        sample_values();
    endtask


    // Function: enable_coverage
    // Build coverage object if it doesn't already exist.
    function void enable_coverage(uvm_reg_cvr_t models, bit cg_per_instance=0);
        if (cg_per_instance) begin
            if (cg == null) begin
                //$info("Creating instance coverage object: %0s", {this.get_full_name(), ".cg"});
                cg = p5_priority_index_reg_cover::type_id::create({this.get_full_name(), ".cg"});
            end
        end else begin
            //$info("Creating singleton coverage object: %0s", {this.get_full_name(), ".cg"});
            cg_all = p5_priority_index_reg_cover::get();
        end
        this.add_coverage(models);
    endfunction


    // Function: sample_values
    // Called in post-actions
    virtual function void sample_values();
        // Sample only if coverage object has been created
        if(cg != null) begin
            cg.sample(this, is_read);
        end
        if (cg_all != null) begin
            cg_all.sample(this, is_read);
        end
    endfunction


    // Function: sample
    // Sample the raw transaction
    //function void sample(uvm_reg_data_t data, uvm_reg_data_t byte_en, bit is_read, uvm_reg_map map);


    // Function: has_params
    function int unsigned has_params();
        has_params = 0;
        has_params += 0;
    endfunction

    // Function: fields2string
    // Stringify fields.
    virtual function string fields2string();
        string s="";
        $swrite(s, "%0s\n%24s=0x%0h", s, if_action_index.get_name, if_action_index.value);
        $swrite(s, "%0s\n%24s=0x%0h", s, cpu_action_index.get_name, cpu_action_index.value);
        $swrite(s, "%0s\n%24s=0x%0h", s, mon1_action_index.get_name, mon1_action_index.value);
        $swrite(s, "%0s\n%24s=0x%0h", s, mon2_action_index.get_name, mon2_action_index.value);
        return s;
    endfunction

endclass


// Class: p5_priority_index_reg_cover
// Register coverage object.
class p5_priority_index_reg_cover extends uvm_object;

    static local p5_priority_index_reg_cover m_inst;

    // Variable: r
    // Handle to register to sample
    p5_priority_index_reg r;

    covergroup cg with function sample(bit is_read);
        option.per_instance = 1;
        type_option.merge_instances = 1;
        if_action_index_wr: coverpoint r.if_action_index.value iff (!is_read) { bins bin[16] = {[0:$]}; }
        if_action_index_rd: coverpoint r.if_action_index.value iff  (is_read) { bins bin[16] = {[0:$]}; }
        cpu_action_index_wr: coverpoint r.cpu_action_index.value iff (!is_read) { bins bin[16] = {[0:$]}; }
        cpu_action_index_rd: coverpoint r.cpu_action_index.value iff  (is_read) { bins bin[16] = {[0:$]}; }
        mon1_action_index_wr: coverpoint r.mon1_action_index.value iff (!is_read);
        mon1_action_index_rd: coverpoint r.mon1_action_index.value iff  (is_read);
        mon2_action_index_wr: coverpoint r.mon2_action_index.value iff (!is_read);
        mon2_action_index_rd: coverpoint r.mon2_action_index.value iff  (is_read);
    endgroup

    `uvm_object_utils(rule_action_mapping_nni10g_reg_pkg::p5_priority_index_reg_cover)

    // Constructor: new
    // Note that to be truly singleton, the constructor should be protected.
    /*protected*/ function new(string name="p5_priority_index_reg_cover");
        super.new(name);
        cg = new(/*name*/);
    endfunction


    // Function: set_name
    // Override function to set name of covergroup.
    virtual function void set_name(string name);
        super.set_name(name);
        cg.option.name = name;
    endfunction


    // Function: get
    // Get the coverage object singleton.
    static function p5_priority_index_reg_cover get();
        if (m_inst == null) begin
            m_inst = p5_priority_index_reg_cover::type_id::create("cg");
        end
        return m_inst;
    endfunction


    // Function: sample
    // Sample the register for coverage.
    virtual function void sample(p5_priority_index_reg _r, bit is_read);
        r = _r;
        cg.sample(is_read);
    endfunction

endclass





// Class: rule_action_mapping_nni10g_reg_block
// Register Block .rule_action_mapping_nni10g: 
class rule_action_mapping_nni10g_reg_block extends uvm_reg_block;

    // Validate register width
    local static bit valid_reg_data_width = check_data_width(`UVM_REG_DATA_WIDTH);

    rand p5_priority_index_reg priority_index[];

    // Variable: params
    // Parameter key/value lookup.
    static protected acd_reg_param_cfg m_params;

    // Variable: cg_per_instance
    // Assert to construct all sub-block and register covergroups per instance rather than singleton
    protected bit cg_per_instance;

    `uvm_object_utils(rule_action_mapping_nni10g_reg_pkg::rule_action_mapping_nni10g_reg_block)

    // Constructor: new
    function new(string name = "rule_action_mapping_nni10g_reg_block");
        super.new(name, UVM_NO_COVERAGE);
    endfunction


    // Function: build
    virtual function void build();
        if ((m_params == null) && (0 > 0))
            if (!uvm_config_db#(acd_reg_param_cfg)::get(null, get_full_name(), "cfg", m_params))
                `uvm_fatal("CFGERR", {get_full_name(), " failed to get configuration for parameters."})

        priority_index = new[4096];

        foreach(priority_index[m]) begin
            priority_index[m] = p5_priority_index_reg::type_id::create($sformatf("priority_index[%0d]",m), , get_full_name());
        end

        foreach(priority_index[m]) begin
            priority_index[m].configure(this);
        end

        foreach(priority_index[m]) begin
            priority_index[m].build();
        end

        // define default map
        default_map = create_map("rule_action_mapping_nni10g_default_map", 'h0, `UVM_REG_DATA_WIDTH/8, UVM_NO_ENDIAN, 0);
        foreach(priority_index[m]) begin
            this.default_map.add_reg(this.priority_index[m], 'h0 + m, "RW");
        end

        // Recursively lock register model and build the address map to enable
        // uvm_reg_map::get_reg_by_offset() and uvm_reg_map::get_mem_by_offset() methods.
        // It is impossible to unlock a model.
        lock_model();
    endfunction


     // Function: set_per_instance_coverage
     // Enable or disable instance coverage, otherwise singleton coverage.
     virtual function void set_per_instance_coverage(bit per_inst, uvm_hier_e hier=UVM_HIER);
         this.cg_per_instance = per_inst;

        // Use UVM_CVR_ALL for hierarchical enabling.
        if(hier == UVM_HIER) begin
        end
     endfunction


    // Function: set_coverage
    // Override base function to create covergroups for all registers in this block.
    //
    // In order to enable hierarchical creation, use UVM_CVR_ALL.
    virtual function uvm_reg_cvr_t set_coverage(uvm_reg_cvr_t is_on);
        //void'(uvm_config_db#(bit)::get(null, get_full_name(), "cg_per_instance", cg_per_instance));
        set_coverage = super.set_coverage(is_on);
        foreach(priority_index[m]) begin
            priority_index[m].enable_coverage(is_on, this.cg_per_instance);
        end
        // Use UVM_CVR_ALL for hierarchical enabling.
        if(is_on == UVM_CVR_ALL) begin
        end
        return set_coverage;
    endfunction


    // Function: fields2string
    // Stringify.
    virtual function string convert2string();
        string s = "";
        uvm_reg regs[$];
        uvm_reg_field fields[$];

        get_registers(regs, UVM_HIER);
        $swrite(s, "\nUVM_REG_BLOCK::%0s (%0d registers)\n", get_name, regs.size());
        foreach (regs[m]) begin
            $swrite(s, "%0s    %0s=0x%16h\n", s, regs[m].get_full_name, regs[m].get());
            // Getting the fields is optional might be too verbose
            //fields.delete();
            //regs[m].get_fields(fields);
            //foreach (fields[n]) begin
                //$swrite(s, "%0s        %0s=0x%0h\n", s, fields[n].get_full_name, fields[n].value);
            //end
        end
        return s;
    endfunction


    // Function: regs2update
    // Stringifying only regmodel registers that need updating. Useful after randomization.
    virtual function string regs2update();
        string s = "";
        uvm_reg regs[$];
        uvm_reg_field fields[$];

        get_registers(regs, UVM_HIER);
        $swrite(s, "\nRegisters requiring update in UVM_REG_BLOCK::%0s\n", get_name);
        foreach (regs[m]) begin
            if (regs[m].needs_update()) begin
                $swrite(s, "%0s    %0s=0x%16h\n", s, regs[m].get_full_name, regs[m].get());
                // Getting the fields is optional might be too verbose
                fields.delete();
                regs[m].get_fields(fields);
                foreach (fields[n]) begin
                    $swrite(s, "%0s        %0s=0x%0h\n", s, fields[n].get_full_name, fields[n].value);
                end
            end
        end
        return s;
    endfunction

endclass

endpackage